class sig_agent_cfg extends hdv_agent_cfg;
  virtual sig_if vif;
  `uvm_object_utils(sig_agent_cfg)

  `uvm_object_new
endclass
