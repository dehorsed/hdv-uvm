package sig_pkg;
  import uvm_pkg::*;
  import hdv_pkg::*;
  `include "sig_agent_cfg.svh"
  `include "sig_seq_item.svh"
  `include "sig_sequencer.svh"
  `include "sig_sequence.svh"
  `include "sig_driver.svh"
  `include "sig_monitor.svh"
  `include "sig_agent.svh"
  `include "sig_scoreboard.svh"
  `include "sig_env.svh"
  `include "sig_test.svh"
endpackage : sig_pkg
