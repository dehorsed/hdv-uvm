class sig_agent extends hdv_pkg::hdv_agent#(sig_agent_cfg, sig_driver, sig_sequencer, sig_monitor, hdv_agent_cov);
  `uvm_component_utils(sig_agent)

  `uvm_component_new
endclass
