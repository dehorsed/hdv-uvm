class sig_sequencer extends hdv_sequencer #(sig_seq_item);
  `uvm_component_utils(sig_sequencer)

  `uvm_component_new

endclass
